----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:25:59 12/01/2018 
-- Design Name: 
-- Module Name:    vga_calc - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
use work.utils.all;

entity vga_calc is
	PORT (
        clk_50, rst: IN STD_LOGIC;
        vga_control_signal: in vga_control;
        data_in: in std_logic_vector(15 downto 0);
        h_sync, v_sync: OUT STD_LOGIC;  --horiztonal, vertical sync pulse
	    r, g, b: out STD_LOGIC_VECTOR(2 downto 0)
	);
end vga_calc;

architecture Behavioral of vga_calc is
	component vga640480 is
		port(
			reset       :         in  STD_LOGIC;
			clk_0       :         in  STD_LOGIC; --50Mʱ������
			hs,vs       :         out STD_LOGIC; --��ͬ������ͬ���ź�
			vector_x_out   :   out std_LOGIC_VECTOR(9 downto 0);  --ɨ��λ�õĺ�����
			vector_y_out :     out std_LOGIC_vector(8 downto 0);  --ɨ��λ�õ�������
			clk25 : out std_logic;  --25Mʱ�����
			q : in std_logic_vector(9 downto 0);
			r,g,b : out std_logic_vector(2 downto 0)
		);
	end component vga640480;
	
	component checkout_pixel is
		port(
			clk: in std_logic;
			disp_data: in std_logic_vector(6 downto 0);
			left_up_point: in point;
			col: in integer;
			row: in integer;
			is_on: out std_logic
		);
	end component checkout_pixel;
	
	signal s_x: std_logic_vector(9 downto 0);
	signal s_y: std_logic_vector(8 downto 0);
	signal clk_25:std_logic;
	signal q_vga: std_logic_vector(9 downto 0);
	
	constant hpStart_x:std_LOGIC_vector(9 downto 0) := "1000111010";
   constant hpEnd_x:std_LOGIC_vector(9 downto 0) := "1001101100";
   constant hpStart_y:std_LOGIC_vector(8 downto 0) := "000010100";
   constant hpEnd_y:std_logic_vector(8 downto 0) := "000011110";
	
	constant FONT_WIDTH: integer:=8;
	constant FONT_HEIGHT: integer:=16;
	 
	signal HpOk: std_logic;		--TODO delete this test
	
	signal disp_data: std_logic_vector(6 downto 0);
	signal left_up_point: point:=(0, 0);
	signal pixel_row, pixel_col : integer;
	signal is_on: std_logic:='0';
	
	signal vga_r, vga_g, vga_b: std_logic_vector(2 downto 0);

	subtype ascii_vec is std_logic_vector(6 downto 0);
	type ascii_vec_array is array(integer range<>) of ascii_vec;
	subtype ascii_col is ascii_vec_array(0 to 79);
	type ascii_col_array is array(integer range<>) of ascii_col;
	subtype ascii_matrix is ascii_col_array(0 to 29);
	
	signal mem: ascii_matrix := (others => (others => (others => '0')));
	
	shared variable cursor_row, cursor_col : integer := 0;
begin
	vga_640480: vga640480
	port map(
		reset => rst,
		clk_0 => clk_50,
		hs => h_sync,
		vs => v_sync,
		vector_x_out => s_x,
		vector_y_out => s_y,
		clk25 => clk_25,
		q => q_vga,
		r => vga_r,
		g => vga_g,
		b => vga_b
	);
	
	check_out_pixel_entity: checkout_pixel
	port map(
		clk => clk_50,
		disp_data => disp_data,
		left_up_point => left_up_point,
		col => pixel_col,
		row => pixel_row,
		is_on => is_on
	);
	
	-------------------------------------------------------------------------
	process(clk_50, s_x, s_y)  --calc pixel col and row
	begin
		if rising_edge(clk_50) then
			pixel_col <= to_integer(unsigned(s_x));
			pixel_row <= to_integer(unsigned(s_y));
		end if;
	end process;
	
	process(clk_50)
	begin
		if rst = '1' then
			cursor_row := 1;
			cursor_col := 0;
			mem <= (others => (others => (others => '0')));
			mem(0)(0) <= std_logic_vector(to_unsigned(character'pos('F'), 7));
			mem(0)(1) <= std_logic_vector(to_unsigned(character'pos('U'), 7));
			mem(0)(2) <= std_logic_vector(to_unsigned(character'pos('C'), 7));
			mem(0)(3) <= std_logic_vector(to_unsigned(character'pos('K'), 7));
		elsif rising_edge(clk_50) then
			case data_in(6 downto 0) is
				when "0001101" => -- Enter
					 cursor_row := cursor_row + 1;
					 cursor_col := 0;
				when "0001000" => -- Backspace
					 mem(cursor_row)(cursor_col) <= (others => '0');
					 cursor_col := cursor_col - 1;
				when others =>
					 mem(cursor_row)(cursor_col) <= data_in(6 downto 0);
					 cursor_col := cursor_col + 1;
					 if cursor_col = 80 then
						  cursor_row := cursor_row + 1;
						  cursor_col := 0;
					 end if;
			end case;
		end if;
	end process;
	
	process(clk_50)
	begin
		if rising_edge(clk_50) then
			left_up_point <= (((pixel_col / FONT_WIDTH) * FONT_WIDTH), ((pixel_row / FONT_HEIGHT) * FONT_HEIGHT));
			if 0 <= pixel_row and pixel_row < 30 * FONT_HEIGHT and 0 <= pixel_col and pixel_col < 80 * FONT_WIDTH then
				disp_data <= mem(pixel_row / FONT_HEIGHT)(pixel_col / FONT_WIDTH);
			else
				disp_data <= "0000000";
			end if;
		end if;
	end process;
	
	
	process(clk_50, is_on)
	begin
		if rising_edge(clk_50) then
			if is_on = '1' then
				q_vga <= "0111111111";
			else
				q_vga <= "0000000000";
			end if;
		end if;
	end process;
	
	process(clk_50, vga_r, vga_b, vga_g)
	begin
		if rising_edge(clk_50) then
			r <= vga_r;
			g <= vga_g;
			b <= vga_b;
		end if;
	end process;
	
	
--	process(clk_50)		--TODO delete this 
--	begin
--		if(s_x >= hpStart_x and s_x <= hpEnd_x and s_y >= hpStart_y and s_y <= hpEnd_y) then
--        if(CONV_INTEGER(s_x - hpStart_x) * 100 <= 100 * 50) then  --������״
--            HpOK <= '1';
--        else
--            HpOK <= '0';
--        end if;
--		else
--        HpOK <= '0';
--		end if;
--	end process;
--	
--	process(clk_25, rst)		--TODO delete this
--	begin
--		if clk_25'event and clk_25 = '1' then
--			if (hpOk = '1') then
--				q_vga <= "0111000000";
--			else
--				q_vga <= "0111111111";
--			end if;
--		end if;
--	end process;
	
end Behavioral;

